module rs_485
#(parameter start_bit = 0, parameter stop_bit = 1)
(
input clk,
input in_data,
output out_strob,
output [7:0] out_data
);



endmodule